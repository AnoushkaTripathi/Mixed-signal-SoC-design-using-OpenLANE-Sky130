magic
tech sky130A
timestamp 1719146560
<< nwell >>
rect 0 291 874 576
<< nmos >>
rect 90 148 110 228
rect 279 148 299 228
rect 665 148 685 228
<< pmos >>
rect 90 360 110 442
rect 279 360 299 442
rect 665 360 685 442
<< ndiff >>
rect 26 211 90 228
rect 26 171 40 211
rect 80 171 90 211
rect 26 148 90 171
rect 110 211 187 228
rect 110 171 120 211
rect 160 171 187 211
rect 110 148 187 171
rect 215 213 279 228
rect 215 173 229 213
rect 269 173 279 213
rect 215 148 279 173
rect 299 213 376 228
rect 299 173 310 213
rect 350 173 376 213
rect 299 148 376 173
rect 602 213 665 228
rect 602 173 616 213
rect 656 173 665 213
rect 602 148 665 173
rect 685 213 763 228
rect 685 173 694 213
rect 734 173 763 213
rect 685 148 763 173
<< pdiff >>
rect 26 423 90 442
rect 26 383 40 423
rect 80 383 90 423
rect 26 360 90 383
rect 110 423 187 442
rect 110 383 121 423
rect 161 383 187 423
rect 110 360 187 383
rect 215 423 279 442
rect 215 383 229 423
rect 269 383 279 423
rect 215 360 279 383
rect 299 423 376 442
rect 299 383 307 423
rect 347 383 376 423
rect 299 360 376 383
rect 602 423 665 442
rect 602 383 616 423
rect 656 383 665 423
rect 602 360 665 383
rect 685 425 763 442
rect 685 385 694 425
rect 734 385 763 425
rect 685 360 763 385
<< ndiffc >>
rect 40 171 80 211
rect 120 171 160 211
rect 229 173 269 213
rect 310 173 350 213
rect 616 173 656 213
rect 694 173 734 213
<< pdiffc >>
rect 40 383 80 423
rect 121 383 161 423
rect 229 383 269 423
rect 307 383 347 423
rect 616 383 656 423
rect 694 385 734 425
<< poly >>
rect 90 450 299 470
rect 90 442 110 450
rect 279 442 299 450
rect 665 442 685 467
rect 90 347 110 360
rect 222 325 257 330
rect 90 322 257 325
rect 90 305 231 322
rect 248 305 257 322
rect 90 294 257 305
rect 90 228 110 294
rect 279 272 299 360
rect 326 339 360 344
rect 665 339 685 360
rect 326 333 685 339
rect 326 316 334 333
rect 351 324 685 333
rect 351 316 360 324
rect 326 308 360 316
rect 245 267 299 272
rect 245 250 254 267
rect 271 250 299 267
rect 245 245 299 250
rect 279 228 299 245
rect 665 228 685 241
rect 90 123 110 148
rect 279 138 299 148
rect 665 138 685 148
rect 279 118 685 138
<< polycont >>
rect 231 305 248 322
rect 334 316 351 333
rect 254 250 271 267
<< locali >>
rect 0 535 15 553
rect 33 535 64 553
rect 82 535 113 553
rect 131 535 162 553
rect 180 535 211 553
rect 229 535 260 553
rect 278 535 309 553
rect 327 535 358 553
rect 376 535 407 553
rect 425 535 456 553
rect 474 535 505 553
rect 523 535 554 553
rect 572 535 603 553
rect 621 535 652 553
rect 670 535 701 553
rect 719 535 750 553
rect 768 535 799 553
rect 817 535 848 553
rect 866 535 874 553
rect 229 440 269 535
rect 28 423 85 440
rect 28 383 40 423
rect 80 383 85 423
rect 28 362 85 383
rect 113 423 185 440
rect 113 383 121 423
rect 161 383 185 423
rect 113 362 185 383
rect 217 423 274 440
rect 217 383 229 423
rect 269 383 274 423
rect 217 362 274 383
rect 302 423 374 440
rect 302 383 307 423
rect 347 383 374 423
rect 302 362 374 383
rect 604 423 661 440
rect 604 383 616 423
rect 656 383 661 423
rect 604 362 661 383
rect 689 425 761 440
rect 689 385 694 425
rect 734 385 761 425
rect 689 362 761 385
rect 40 228 80 362
rect 121 228 160 362
rect 310 345 350 362
rect 247 344 350 345
rect 247 333 360 344
rect 247 330 334 333
rect 222 322 334 330
rect 222 305 231 322
rect 248 316 334 322
rect 351 316 360 333
rect 248 308 360 316
rect 248 305 350 308
rect 222 294 257 305
rect 292 304 350 305
rect 177 259 191 277
rect 209 259 228 277
rect 245 267 280 272
rect 245 250 254 267
rect 271 250 280 267
rect 245 245 280 250
rect 28 211 85 228
rect 28 171 40 211
rect 80 171 85 211
rect 28 150 85 171
rect 113 211 185 228
rect 113 171 120 211
rect 160 171 185 211
rect 203 214 211 225
rect 310 226 350 304
rect 367 259 382 277
rect 400 259 431 277
rect 449 259 480 277
rect 498 259 529 277
rect 547 259 578 277
rect 596 259 599 277
rect 616 226 656 362
rect 694 226 734 362
rect 751 259 766 277
rect 784 259 815 277
rect 833 259 874 277
rect 228 214 274 226
rect 203 213 274 214
rect 203 200 229 213
rect 113 150 185 171
rect 217 173 229 200
rect 269 173 274 213
rect 217 150 274 173
rect 302 213 374 226
rect 302 173 310 213
rect 350 173 374 213
rect 302 150 374 173
rect 604 213 661 226
rect 604 173 616 213
rect 656 173 661 213
rect 604 150 661 173
rect 689 213 761 226
rect 689 173 694 213
rect 734 173 761 213
rect 689 150 761 173
rect 120 119 160 150
rect 616 119 656 150
rect 120 102 656 119
rect 0 -9 15 9
rect 33 -9 64 9
rect 82 -9 113 9
rect 131 -9 162 9
rect 180 -9 211 9
rect 229 -9 260 9
rect 278 -9 309 9
rect 327 -9 358 9
rect 376 -9 407 9
rect 425 -9 456 9
rect 474 -9 505 9
rect 523 -9 554 9
rect 572 -9 603 9
rect 621 -9 652 9
rect 670 -9 701 9
rect 719 -9 750 9
rect 768 -9 799 9
rect 817 -9 848 9
rect 866 -9 872 9
<< viali >>
rect 15 535 33 553
rect 64 535 82 553
rect 113 535 131 553
rect 162 535 180 553
rect 211 535 229 553
rect 260 535 278 553
rect 309 535 327 553
rect 358 535 376 553
rect 407 535 425 553
rect 456 535 474 553
rect 505 535 523 553
rect 554 535 572 553
rect 603 535 621 553
rect 652 535 670 553
rect 701 535 719 553
rect 750 535 768 553
rect 799 535 817 553
rect 848 535 866 553
rect 191 259 209 277
rect 211 214 228 231
rect 382 259 400 277
rect 431 259 449 277
rect 480 259 498 277
rect 529 259 547 277
rect 578 259 596 277
rect 766 259 784 277
rect 815 259 833 277
rect 15 -9 33 9
rect 64 -9 82 9
rect 113 -9 131 9
rect 162 -9 180 9
rect 211 -9 229 9
rect 260 -9 278 9
rect 309 -9 327 9
rect 358 -9 376 9
rect 407 -9 425 9
rect 456 -9 474 9
rect 505 -9 523 9
rect 554 -9 572 9
rect 603 -9 621 9
rect 652 -9 670 9
rect 701 -9 719 9
rect 750 -9 768 9
rect 799 -9 817 9
rect 848 -9 866 9
<< metal1 >>
rect 0 553 874 568
rect 0 535 15 553
rect 33 535 64 553
rect 82 535 113 553
rect 131 535 162 553
rect 180 535 211 553
rect 229 535 260 553
rect 278 535 309 553
rect 327 535 358 553
rect 376 535 407 553
rect 425 535 456 553
rect 474 535 505 553
rect 523 535 554 553
rect 572 535 603 553
rect 621 535 652 553
rect 670 535 701 553
rect 719 535 750 553
rect 768 535 799 553
rect 817 535 848 553
rect 866 535 874 553
rect 0 520 874 535
rect 0 277 874 292
rect 0 259 191 277
rect 209 259 382 277
rect 400 259 431 277
rect 449 259 480 277
rect 498 259 529 277
rect 547 259 578 277
rect 596 259 766 277
rect 784 259 815 277
rect 833 259 874 277
rect 0 244 874 259
rect 203 231 242 244
rect 203 214 211 231
rect 228 225 242 231
rect 228 214 245 225
rect 203 200 245 214
rect 0 9 872 24
rect 0 -9 15 9
rect 33 -9 64 9
rect 82 -9 113 9
rect 131 -9 162 9
rect 180 -9 211 9
rect 229 -9 260 9
rect 278 -9 309 9
rect 327 -9 358 9
rect 376 -9 407 9
rect 425 -9 456 9
rect 474 -9 505 9
rect 523 -9 554 9
rect 572 -9 603 9
rect 621 -9 652 9
rect 670 -9 701 9
rect 719 -9 750 9
rect 768 -9 799 9
rect 817 -9 848 9
rect 866 -9 872 9
rect 0 -24 872 -9
<< labels >>
flabel locali s 59 284 59 284 0 FreeSans 120 0 0 0 I1
port 14 nsew signal input
<< properties >>
string LEFclass CORE
string LEFsite unithdbl LEForigin 0 0
string FIXED_BBOX 0 0 874 544
<< end >>
